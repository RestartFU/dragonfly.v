module main

import server

fn main() {
	mut s := server.new()!
	for {
		mut p, ok := s.accept()
		if !ok {
			return
		}
		p.message("welcome, ${p.name()}")
		mut player_list := []string{}
		for mut pl in s.players() {
			player_list << pl.name()
		}
		println("players online: ${player_list.join(", ")}")
	}
}
